module ram_memory(    
    input reset, 
    input [25:0] data_requested,where_to_write,
    output reg [127:0] data_returned,
    input [127:0] data_to_write,
    input write_to_mem);

    reg [31:0] memory [10485:0]; //han de ser 20 bits per addreces fisiques

    reg [31:0] shifted_adress,shifted_adress_write;
    int k,j;
    always @ (*) begin
        
        if (reset == 1'b1) begin
            /*for (int i=0; i < 1048576; i++) begin
                memory[i] = i;
            end*/
            /*memory[0] <=   32'b000010_00000000010000001000001010;
            memory[1] <=   32'b000000_00000000110011000000000010;
            memory[2] <=   32'b000000_00000110001010010100011000;
            memory[3] <=   32'b000010_00000000000000111000001010;
            memory[4] <=   32'b000010_00000_11111_0000000000000000;
            memory[5] <=   32'b000100_11111_10000_0001_0000_0000_0000; // LD R16 <- 0(R31) 0x1000 //4096
            memory[6] <=   32'b000010_00000000010000001000001010;
            memory[7] <=   32'b000000_00000000110011000000000010;
            memory[8] <=   32'b000000_00000110001010010100011000;
            memory[9] <=   32'b000010_00000000000000111000001010;*/



            memory[0] = 32'b000010_00000_00001_0000_0000_1000_0000; // ADDI R1 <- R0,0x80 //128
            memory[1] = 32'b000010_00000_11111_0000_0000_0000_0000; // ADDI R31 <- R0,0x00 //0
            memory[2] = 32'b000010_00000_00101_0000_0000_0000_0000; // ADDI R5 <- R0,0x00 //0 i
            memory[3] = 32'b000010_00000_00010_0000_0000_0000_0000; // ADDI R2 <- R0,0x00 //0 count
            memory[4] = 32'b000100_00010_00011_0010_0000_0000_0000; // LD R3 <- 0x2000(R2)
            memory[5] = 32'b000000_00011_11111_11111_000_0000_0010; // ADD R31 <- R3,R31
            memory[6] = 32'b000010_00000_00010_0000_0000_0000_0100; // ADDI R2 <- R0,0x04 //4 ++count
            memory[7] = 32'b000010_00000_00101_0000_0000_0000_0001; // ADDI R5 <- R0,0x01 //1 ++count
            memory[8] = 32'b000000_00101_00110_00101_00000001000; // COMPLT R6 <- R5, R1
            memory[9] = 32'b001001_00110_00000_000_0000_0000_000; // BEQ R6,R0, 0x000
            
            //sore_buffer + data_cache
            /*memory[0] <=   32'b00000000000000000000000000000000;
            memory[1] <=   32'b00000000000000000000000000000001;
            memory[2] <=   32'b00000000000000000000000000000010;
            memory[3] <=   32'b00000000000000000000000000000110;
            memory[4] <=   32'b00000000000000000000000000000100;
            memory[5] <=   32'b00000000000000000000000000000101;
            memory[6] <=   32'b00000000000000000000000000000110;
            memory[7] <=   32'b00000000000000000000000000000111;
            memory[8] <=   32'b00000000000000000000000000001000;
            memory[9] <=   32'b00000000000000000000000000001001;
            memory[10] <=  32'b00000000000000000000000000001010;
            memory[11] <=  32'b00000000000000000000000000001011;
            memory[12] <=  32'b00000000000000000000000000001100;
            memory[13] <=  32'b00000000000000000000000000001101;
            memory[14] <=  32'b00000000000000000000000000001110;
            memory[15] <=  32'b00000000000000000000000000001111;
            memory[16] <=  32'b00000000000000000000000000010000;
            memory[17] <=  32'b00000000000000000000000000010001;
            memory[18] <=  32'b00000000000000000000000000010010;
            memory[19] <=  32'b00000000000000000000000000010011;
            memory[20] <=  32'b00000000000000000000000000010100;
            memory[21] <=  32'b00000000000000000000000000010101;
            memory[22] <=  32'b00000000000000000000000000010110;
            memory[23] <=  32'b00000000000000000000000000010111;
            memory[24] <=  32'b00000000000000000000000000011000;
            memory[25] <=  32'b00000000000000000000000000011001;
            memory[26] <=  32'b00000000000000000000000000011010;
            memory[27] <=  32'b00000000000000000000000000011011;
            memory[28] <=  32'b00000000000000000000000000011100;
            memory[29] <=  32'b00000000000000000000000000011101;
            memory[30] <=  32'b00000000000000000000000000011110;
            memory[31] <=  32'b00000000000000000000000000011111;
            memory[32] <=  32'b00000000000000000000000000100001;
            memory[33] <=  32'b00000000000000000000000000100010;
            memory[34] <=  32'b00000000000000000000000000100011;
            memory[35] <=  32'b00000000000000000000000000100100;
            memory[36] <=  32'b00000000000000000000000000100101;
            memory[37] <=  32'b00000000000000000000000000100110;
            memory[38] <=  32'b00000000000000000000000000100111;
            memory[39] <=  32'b00000000000000000000000000101000;
            memory[40] <=  32'b00000000000000000000000000101001;
            memory[41] <=  32'b00000000000000000000000000101010;
            memory[42] <=  32'b00000000000000000000000000101011;
            memory[43] <=  32'b00000000000000000000000000101100;
            memory[44] <=  32'b00000000000000000000000000101101;
            memory[45] <=  32'b00000000000000000000000000101110;
            memory[46] <=  32'b00000000000000000000000000101111;
            memory[47] <=  32'b00000000000000000000000000110000;
            memory[48] <=  32'b00000000000000000000000000110001;
            memory[49] <=  32'b00000000000000000000000000110010;
            memory[50] <=  32'b00000000000000000000000000110011;
            memory[51] <=  32'b00000000000000000000000000110100;*/
            memory[4096] =   32'b000000_00000_00000_0000_0000_0000_0000;
            memory[8192] =   32'b000000_00000_00000_0000_0000_0000_0000;
            memory[8193] =   32'b000000_00000_00000_0000_0000_0000_0000;
            memory[8194] =   32'b000000_00000_00000_0000_0000_0000_0000;
            memory[8195] =   32'b000000_00000_00000_0000_0000_0000_0000;
            k = 8192;
            for (int i = 0; i < 128; i++) begin
                j = k + i;
                memory[j] = i;
            end

        end
        
        else begin
            shifted_adress = data_requested << 2;
            data_returned = {memory[shifted_adress + 3], memory[shifted_adress + 2], memory[shifted_adress + 1], memory[shifted_adress]};
            if (write_to_mem == 1'b1) begin
                shifted_adress_write = where_to_write << 2;
                {memory[shifted_adress_write + 3], memory[shifted_adress_write + 2], memory[shifted_adress_write + 1], memory[shifted_adress_write]} = data_to_write;
            end
        end

    end

endmodule // insttructionMem





/*

        memory[0] = 000010_00000_00001_0000_0000_1000_0000; // ADDI R1 <- R0,0x80 //128
        memory[1] = 000010_00000_11111_0000_0000_0000_0000; // ADDI R31 <- R0,0x00 //0
        memory[2] = 000010_00000_00101_0000_0000_0000_0000; // ADDI R5 <- R0,0x00 //0 i
        memory[3] = 000010_00000_00010_0000_0000_0000_0000; // ADDI R2 <- R0,0x00 //0 count
        memory[4] = 000100_00010_00011_0010_0000_0000_0000; // LD R3 <- 0x2000(R2)
        memory[5] = 000000_00011_11111_11111_0000_0000_0010; // ADD R31 <- R3,R31
        memory[6] = 000010_00000_00010_0000_0000_0000_0100; // ADDI R2 <- R0,0x04 //4 ++count
        memory[7] = 000010_00000_00010_0000_0000_0000_0001; // ADDI R2 <- R0,0x01 //1 ++count
        memory[8] = 000000_00101_00110_00101_000000001000; // COMPLT R6 <- R5, R1
        memory[9] = 001001_00110_00000_000_0000_0000_0000; // BEQ R6,R0, 0x000


*/